40
8
30
9750
