15
-3
45
15000
