50
15
-3
45
5000
