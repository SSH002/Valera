0
-3
100
28750
